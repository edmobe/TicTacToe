library verilog;
use verilog.vl_types.all;
entity testbench_Top is
end testbench_Top;
