library verilog;
use verilog.vl_types.all;
entity testbench_Sprite_Controller is
end testbench_Sprite_Controller;
