library verilog;
use verilog.vl_types.all;
entity testbench_Sram is
end testbench_Sram;
