`timescale 1ns / 1ps
// Counter based
module clock_divider #(parameter div_value = 1) (
	input logic clk, // 100 MHz
	output logic divided_clk = 0 // 25 MHz
);

	// Division value = 100 MHz / (2 * desired frequency) - 1
	// Counter
	integer counter_value = 0; // 32 bit wide bus

	always @ (posedge clk)
	begin
		// Keep counting until division
		if (counter_value == div_value)
			counter_value = 0;
		else
			counter_value = counter_value + 1;
	end

	// Divide clock
	always @ (posedge clk)
	begin
		// Keep counting until division
		if (counter_value == div_value)
			divided_clk = ~divided_clk;
		else
			divided_clk = divided_clk;
	end
endmodule
