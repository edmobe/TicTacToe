library verilog;
use verilog.vl_types.all;
entity testbench_TicTacToe is
end testbench_TicTacToe;
