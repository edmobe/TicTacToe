library verilog;
use verilog.vl_types.all;
entity testbench_Video_Controller is
end testbench_Video_Controller;
